adress
ambulans
antenn
backar
bakar
biljett
blåklocka
byte
dagboken
daggmask
docka
dockor
dricka
dörrmatta
ficka
fjäril
flyta
flytta
färggrann
färggrant
glas
glasögon
granbarren
grovt
gryta
grytor
gräddglass
gul
gulare
gulast
halvt
handduk
håla
högt
kamma
karott
kasta
kastade
kastat
krama
kulor
lilla
limpa
limpor
madrass
manet
maskros
mata
matta
mysigt
måne
mätta
noggrann
noggrant
nummer
numret
nötter
parkett
present
pupill
påminde
påminna
påmint
racket
ridstövlar
rosett
ryker
servett
sillar
skalen
skolbuss
skutta
smörgås
snabbt
solros
sommar
somrar
spela
spelade
spelat
spenat
staket
styggt
syren
tallar
tallen
tennis
tofsar
trappa
tändsticka
villa
väggklocka
äggkopp
ögon

banan
biljett
bock
bok
boll
brevet
bromsat
brun
brunn
bullar
bus
buss
citron
dag
dam
damm
dörr
fiskar
flagga
flaggor
flicka
flitig
flyta
gardin
gata
glas
glass
granar
gratis
huset
hög
högg
kakor
kapten
katt
klocka
klockor
klubba
klubbor
knapp
knuffat
komet
kopp
krock
krona
kronor
kropp
lamm
lapp
listig
lock
lok
lykta
lyktor
lönn
lös
löss
lövet
maten
melon
myra
myror
nyckel
näbb
och
också
pojke
raket
repet
rida
rider
ryka
ryker
rönn
sitta
sitter
skalar
skola
sladd
spann
stopp
straff
sågar
tabell
taggig
taket
trollet
trumpet
tulpan
tupp
tältar
vispar
vulkan
vägg
ägg
ägget

arm
bok
brud
bur
båt
dag
dagg
fat
fest
fisk
fot
glas
glass
gräs
gröt
hall
han
hett
hon
hål
häl
hök
jal
kan
knyst
ko
kor
kram
kräm
kör
lag
lätt
lök
mest
min
mus
mås
nål
nöt
par
press
rygg
rök
skål
slöjd
sol
stol
stress
sår
sås
söt
tak
tal
tall
trygg
tråd
träd
tub
tyst
tåg
tät
ur
vas
vass
våg
väg
vän
väst
ål
ärm
